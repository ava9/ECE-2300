library verilog;
use verilog.vl_types.all;
entity lab4_test is
end lab4_test;

library verilog;
use verilog.vl_types.all;
entity lab3_test is
end lab3_test;
